library verilog;
use verilog.vl_types.all;
entity Odev_1_vlg_check_tst is
    port(
        BUS_1           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Odev_1_vlg_check_tst;
