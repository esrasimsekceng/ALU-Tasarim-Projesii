library verilog;
use verilog.vl_types.all;
entity Odev_1_vlg_vec_tst is
end Odev_1_vlg_vec_tst;
